*** SPICE deck for cell GDI_Comparator{sch} from library GDI
*** Created on Tue May 21, 2024 23:46:41
*** Last revised on Thu Jun 06, 2024 00:29:52
*** Written on Thu Jun 06, 2024 00:42:55 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT GDI_tech__2And FROM CELL GDI_tech:2And{sch}
.SUBCKT GDI_tech__2And A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 out A B gnd NMOS L=45nm W=4.5U
Mpmos-4@0 gnd A out vdd PMOS L=45nm W=9U
.ENDS GDI_tech__2And

*** SUBCIRCUIT GDI_tech__2XOR FROM CELL GDI_tech:2XOR{sch}
.SUBCKT GDI_tech__2XOR A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@21 B gnd gnd NMOS L=45nm W=90nm
Mnmos-4@1 out A net@21 gnd NMOS L=45nm W=90nm
Mpmos-4@0 vdd B net@21 vdd PMOS L=45nm W=180nm
Mpmos-4@1 B A out vdd PMOS L=45nm W=180nm
.ENDS GDI_tech__2XOR

*** SUBCIRCUIT GDI_tech__3And FROM CELL GDI_tech:3And{sch}
.SUBCKT GDI_tech__3And A B C out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@37 A B gnd NMOS L=45nm W=90nm
Mnmos-4@1 out C net@37 gnd NMOS L=45nm W=135nm
Mpmos-4@0 gnd A net@37 vdd PMOS L=45nm W=180nm
Mpmos-4@1 gnd C out vdd PMOS L=45nm W=270nm
.ENDS GDI_tech__3And

*** SUBCIRCUIT GDI_tech__4And FROM CELL GDI_tech:4And{sch}
.SUBCKT GDI_tech__4And A B C D out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@28 A B gnd NMOS L=45nm W=90nm
Mnmos-4@1 net@52 C net@28 gnd NMOS L=45nm W=135nm
Mnmos-4@2 out net@52 D gnd NMOS L=45nm W=200nm
Mpmos-4@0 gnd A net@28 vdd PMOS L=45nm W=180nm
Mpmos-4@1 gnd C net@52 vdd PMOS L=45nm W=270nm
Mpmos-4@2 gnd net@52 out vdd PMOS L=45nm W=400nm
.ENDS GDI_tech__4And

*** SUBCIRCUIT GDI_tech__5OR FROM CELL GDI_tech:5OR{sch}
.SUBCKT GDI_tech__5OR A B C D E out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@108 A vdd gnd NMOS L=45nm W=90nm
Mnmos-4@1 net@118 C vdd gnd NMOS L=45nm W=90nm
Mnmos-4@2 net@131 D vdd gnd NMOS L=45nm W=90nm
Mnmos-4@3 out E vdd gnd NMOS L=45nm W=90nm
Mpmos-4@0 B A net@108 vdd PMOS L=45nm W=180nm
Mpmos-4@1 net@108 C net@118 vdd PMOS L=45nm W=180nm
Mpmos-4@2 net@118 D net@131 vdd PMOS L=45nm W=180nm
Mpmos-4@3 net@131 E out vdd PMOS L=45nm W=180nm
.ENDS GDI_tech__5OR

*** SUBCIRCUIT GDI_tech__And-5 FROM CELL GDI_tech:And-5{sch}
.SUBCKT GDI_tech__And-5 A B C D E out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 net@375 A B gnd NMOS L=45nm W=90nm
Mnmos-4@1 net@380 C net@375 gnd NMOS L=45nm W=135nm
Mnmos-4@2 net@385 D net@380 gnd NMOS L=45nm W=200nm
Mnmos-4@3 out E net@385 gnd NMOS L=45nm W=300nm
Mpmos-4@0 gnd A net@375 vdd PMOS L=45nm W=180nm
Mpmos-4@1 gnd C net@380 vdd PMOS L=45nm W=270nm
Mpmos-4@2 gnd D net@385 vdd PMOS L=45nm W=400nm
Mpmos-4@3 gnd E out vdd PMOS L=45nm W=600nm
.ENDS GDI_tech__And-5

*** SUBCIRCUIT GDI_tech__inverter FROM CELL GDI_tech:inverter{sch}
.SUBCKT GDI_tech__inverter A out
** GLOBAL gnd
** GLOBAL vdd
Mnmos-4@0 out A gnd gnd NMOS L=45nm W=4.5U
Mpmos-4@0 vdd A out vdd PMOS L=45nm W=9U
.ENDS GDI_tech__inverter

.global gnd vdd

*** TOP LEVEL CELL: GDI_Comparator{sch}
X_2And@4 A3 net@549 net@795 GDI_tech__2And
X_2And@5 net@550 net@663 net@789 GDI_tech__2And
X_2And@6 net@554 B3 net@699 GDI_tech__2And
X_2And@7 net@663 net@667 net@673 GDI_tech__2And
X_2XOR@5 A3 B3 A2 GDI_tech__2XOR
X_2XOR@6 A2 B2 net@541 GDI_tech__2XOR
X_2XOR@7 net@550 B1 net@539 GDI_tech__2XOR
X_2XOR@8 A0 B0 net@540 GDI_tech__2XOR
X_3And@3 net@744 _3And@3_B A2 net@798 GDI_tech__3And
X_3And@4 net@569 B2 A2 net@704 GDI_tech__3And
X_4And@2 net@541 A2 A1 net@788 net@802 GDI_tech__4And
X_4And@3 net@541 A2 net@606 B0 net@707 GDI_tech__4And
X_5OR@2 net@795 net@798 net@802 net@806 net@809 G0 GDI_tech__5OR
X_5OR@3 net@699 net@704 net@707 net@713 net@715 L0 GDI_tech__5OR
XAnd-5@5 A2 net@541 net@539 A0 net@712 net@806 GDI_tech__And-5
XAnd-5@6 A2 net@541 net@539 net@540 net@789 net@809 GDI_tech__And-5
XAnd-5@7 A2 net@541 net@539 net@540 Ei E0 GDI_tech__And-5
XAnd-5@8 A2 net@541 net@539 net@638 B0 net@713 GDI_tech__And-5
XAnd-5@9 net@540 net@673 A2 net@541 net@539 net@715 GDI_tech__And-5
Xinverter@13 B0 net@712 GDI_tech__inverter
Xinverter@14 A0 net@638 GDI_tech__inverter
Xinverter@15 B1 net@788 GDI_tech__inverter
Xinverter@16 A1 net@606 GDI_tech__inverter
Xinverter@17 B2 net@744 GDI_tech__inverter
Xinverter@18 A2 net@569 GDI_tech__inverter
Xinverter@19 B3 net@549 GDI_tech__inverter
Xinverter@20 A3 net@554 GDI_tech__inverter
Xinverter@21 Ei net@663 GDI_tech__inverter
Xinverter@22 Li net@550 GDI_tech__inverter
Xinverter@23 Gi net@667 GDI_tech__inverter

* Spice Code nodes in cell cell 'GDI_Comparator{sch}'
V3 Gi 0 DC 1.8 PULSE 0 1.8 0 0 1ps 1ps 100ns 200ns
V4 Ei 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 50ns 100ns
V6 Li 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 25ns 50ns
V7 A3 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 30ns 70ns
V8 A2 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 40ns 90ns
V9 A1 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 20ns 50ns
V10 A0 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 30ns 60ns
V11 B3 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 20ns 40ns
V12 B2 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 20ns 80ns
V13 B1 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 30ns 70ns
V14 B0 0 DC 1.8 PULSE 1.8 0 0 1ps 1ps 40ns 80ns
.tran 1ps 200ns
V0 VDD 0 DC 1.8
.include C:\Users\a-ahm\Desktop\C5_models.txt
.END
